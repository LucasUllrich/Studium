----------------------------------------------------------------------------
-- Title      : VGA Control
-- Project    : VGA Controller
----------------------------------------------------------------------------
-- File       : vga_control_rtl_cfg.vhd
-- Author     : Lucas Ullrich
-- Company    : FH Technikum Wien, BEL
-- Last update: <date>
-- Platform   : ModelSim, Xilinx Vivado, Basys3
----------------------------------------------------------------------------
-- Description: <What is this code for?>
----------------------------------------------------------------------------
-- Revisions  :
-- Date         Version       Author          Description
-- <date>       <nr.>         Lucas Ullrich   <changes done>
----------------------------------------------------------------------------

configuration vga_control_rtl_cfg of vga_control is
  for rtl
  end for;
end vga_control_rtl_cfg;
