----------------------------------------------------------------------------
-- Title      : Prescaler
-- Project    : VGA Controller
----------------------------------------------------------------------------
-- File       : prescaler.vhd
-- Author     : Lucas Ullrich
-- Company    : FH Technikum Wien, BEL
-- Last update: <date>
-- Platform   : ModelSim, Xilinx Vivado, Basys3
----------------------------------------------------------------------------
-- Description: <What is this code for?>
----------------------------------------------------------------------------
-- Revisions  :
-- Date         Version       Author          Description
-- <date>       <nr.>         Lucas Ullrich   <changes done>
----------------------------------------------------------------------------

configuration prescaler_rtl_cfg of prescaler is
  for rtl
  end for;
end prescaler_rtl_cfg;
