----------------------------------------------------------------------------
-- Title      : Picture Memory Controller
-- Project    : VGA Controller
----------------------------------------------------------------------------
-- File       : tb_mem_ctrl_pic_sim_cfg.vhd
-- Author     : Lucas Ullrich
-- Company    : FH Technikum Wien, BEL
-- Last update: <date>
-- Platform   : ModelSim, Xilinx Vivado, Basys3
----------------------------------------------------------------------------
-- Description: <What is this code for?>
----------------------------------------------------------------------------
-- Revisions  :
-- Date         Version       Author          Description
-- <date>       <nr.>         Lucas Ullrich   <changes done>
----------------------------------------------------------------------------
